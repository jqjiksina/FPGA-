module tb_ddr3(

   );
endmodule